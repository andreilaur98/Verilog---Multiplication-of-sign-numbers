module multiplier(
	input [14:0] x,
	input [14:0] y,
	output[14:0] product
    );
	 
	 reg[3:0] i;
	 reg[7:0] s,d;
	 reg [16:0] A;
	 reg [16:0] S;
	 reg [16:0] P;

	reg signed [7:0] s1,s2,d1,d2,s3,s4,d3,d4,s5,d5;
	reg schimba=0;

always@(*) begin //decodificari
	//cifra din dreapta pt primul nr
	if(x[0]==0 && x[1]==1 && x[2]==1 && x[3]==1 && x[4]==1 && x[5]==1 && x[6]==1)
		s2=8'b00000000;
	if(x[0]==0 && x[1]==0 && x[2]==0 && x[3]==0 && x[4]==1 && x[5]==1 && x[6]==0)
		s2=8'b00000001;
	if(x[0]==1 && x[1]==0 && x[2]==1 && x[3]==1 && x[4]==0 && x[5]==1 && x[6]==1)
		s2=8'b00000010;	
	if(x[0]==1 && x[1]==0 && x[2]==0 && x[3]==1 && x[4]==1 && x[5]==1 && x[6]==1)
		s2=8'b00000011;	
	if(x[0]==1 && x[1]==1 && x[2]==0 && x[3]==0 && x[4]==1 && x[5]==1 && x[6]==0)
		s2=8'b00000100;
	if(x[0]==1 && x[1]==1 && x[2]==0 && x[3]==1 && x[4]==1 && x[5]==0 && x[6]==1)
		s2=8'b00000101;
	if(x[0]==1 && x[1]==1 && x[2]==1 && x[3]==1 && x[4]==1 && x[5]==0 && x[6]==1)
		s2=8'b00000110;
	if(x[0]==0 && x[1]==0 && x[2]==0 && x[3]==0 && x[4]==1 && x[5]==1 && x[6]==1)
		s2=8'b00000111;
	if(x[0]==1 && x[1]==1 && x[2]==1 && x[3]==1 && x[4]==1 && x[5]==1 && x[6]==1)
		s2=8'b00001000;
	if(x[0]==1 && x[1]==1 && x[2]==0 && x[3]==1 && x[4]==1 && x[5]==1 && x[6]==1)
		s2=8'b00001001;
		
	//cifra din stanga pt primul nr
	if(x[7]==0 && x[8]==1 && x[9]==1 && x[10]==1 && x[11]==1 && x[12]==1 && x[13]==1)
		s1=8'b00000000;
	if(x[7]==0 && x[8]==0 && x[9]==0 && x[10]==0 && x[11]==1 && x[12]==1 && x[13]==0)
		s1=8'b00000001;
	if(x[7]==1 && x[8]==0 && x[9]==1 && x[10]==1 && x[11]==0 && x[12]==1 && x[13]==1)
		s1=8'b00000010;	
	if(x[7]==1 && x[8]==0 && x[9]==0 && x[10]==1 && x[11]==1 && x[12]==1 && x[13]==1)
		s1=8'b00000011;	
	if(x[7]==1 && x[8]==1 && x[9]==0 && x[10]==0 && x[11]==1 && x[12]==1 && x[13]==0)
		s1=8'b00000100;
	if(x[7]==1 && x[8]==1 && x[9]==0 && x[10]==1 && x[11]==1 && x[12]==0 && x[13]==1)
		s1=8'b00000101;
	if(x[7]==1 && x[8]==1 && x[9]==1 && x[10]==1 && x[11]==1 && x[12]==0 && x[13]==1)
		s1=8'b00000110;
	if(x[7]==0 && x[8]==0 && x[9]==0 && x[10]==0 && x[11]==1 && x[12]==1 && x[13]==1)
		s1=8'b00000111;
	if(x[7]==1 && x[8]==1 && x[9]==1 && x[10]==1 && x[11]==1 && x[12]==1 && x[13]==1)
		s1=8'b00001000;
	if(x[7]==1 && x[8]==1 && x[9]==0 && x[10]==1 && x[11]==1 && x[12]==1 && x[13]==1)
		s1=8'b00001001;	
		
	//cifra din dreapta pt al 2lea nr
	if(y[0]==0 && y[1]==1 && y[2]==1 && y[3]==1 && y[4]==1 && y[5]==1 && y[6]==1)
		d2=8'b00000000;
	if(y[0]==0 && y[1]==0 && y[2]==0 && y[3]==0 && y[4]==1 && y[5]==1 && y[6]==0)
		d2=8'b00000001;
	if(y[0]==1 && y[1]==0 && y[2]==1 && y[3]==1 && y[4]==0 && y[5]==1 && y[6]==1)
		d2=8'b00000010;	
	if(y[0]==1 && y[1]==0 && y[2]==0 && y[3]==1 && y[4]==1 && y[5]==1 && y[6]==1)
		d2=8'b00000011;	
	if(y[0]==1 && y[1]==1 && y[2]==0 && y[3]==0 && y[4]==1 && y[5]==1 && y[6]==0)
		d2=8'b00000100;
	if(y[0]==1 && y[1]==1 && y[2]==0 && y[3]==1 && y[4]==1 && y[5]==0 && y[6]==1)
		d2=8'b00000101;
	if(y[0]==1 && y[1]==1 && y[2]==1 && y[3]==1 && y[4]==1 && y[5]==0 && y[6]==1)
		d2=8'b00000110;
	if(y[0]==0 && y[1]==0 && y[2]==0 && y[3]==0 && y[4]==1 && y[5]==1 && y[6]==1)
		d2=8'b00000111;
	if(y[0]==1 && y[1]==1 && y[2]==1 && y[3]==1 && y[4]==1 && y[5]==1 && y[6]==1)
		d2=8'b00001000;
	if(y[0]==1 && y[1]==1 && y[2]==0 && y[3]==1 && y[4]==1 && y[5]==1 && y[6]==1)
		d2=8'b00001001;
		
	//cifra din stanga pt al doilea nr
	if(y[7]==0 && y[8]==1 && y[9]==1 && y[10]==1 && y[11]==1 && y[12]==1 && y[13]==1)
		d1=8'b00000000;
	if(y[7]==0 && y[8]==0 && y[9]==0 && y[10]==0 && y[11]==1 && y[12]==1 && y[13]==0)
		d1=8'b00000001;
	if(y[7]==1 && y[8]==0 && y[9]==1 && y[10]==1 && y[11]==0 && y[12]==1 && y[13]==1)
		d1=8'b00000010;	
	if(y[7]==1 && y[8]==0 && y[9]==0 && y[10]==1 && y[11]==1 && y[12]==1 && y[13]==1)
		d1=8'b00000011;	
	if(y[7]==1 && y[8]==1 && y[9]==0 && y[10]==0 && y[11]==1 && y[12]==1 && y[13]==0)
		d1=8'b00000100;
	if(y[7]==1 && y[8]==1 && y[9]==0 && y[10]==1 && y[11]==1 && y[12]==0 && y[13]==1)
		d1=8'b00000101;
	if(y[7]==1 && y[8]==1 && y[9]==1 && y[10]==1 && y[11]==1 && y[12]==0 && y[13]==1)
		d1=8'b00000110;
	if(y[7]==0 && y[8]==0 && y[9]==0 && y[10]==0 && y[11]==1 && y[12]==1 && y[13]==1)
		d1=8'b00000111;
	if(y[7]==1 && y[8]==1 && y[9]==1 && y[10]==1 && y[11]==1 && y[12]==1 && y[13]==1)
		d1=8'b00001000;
	if(y[7]==1 && y[8]==1 && y[9]==0 && y[10]==1 && y[11]==1 && y[12]==1 && y[13]==1)
		d1=8'b00001001;	
	
	// formarea numarului din stanga in binar	
	s3=s1<<3;
	s4=s1<<1;
	s5=s3+s4;
	s=s5+s2;
	
	//formarea numarului din dreapta in binar
	d3=d1<<3;
	d4=d1<<1;
	d5=d3+d4;
	d=d5+d2;
end		


//alg Booth	

always @(*) begin
	if(x[14]==1)
		begin
	A={-s, 9'b000000000};
	S={s, 9'b000000000};
		end
	else 
		begin
	A={s, 9'b000000000};
	S={-s, 9'b000000000};
		end
	
	if(y[14]==1) begin
		P={8'b00000000,-d,1'b0};
	end
		else begin
		P={8'b00000000,d,1'b0};
	end
	
	for(i=0;i<8;i=i+1) begin
	
		case(P[1:0])
	
		2'b00,2'b11:begin
			schimba=P[16];
			P=P>>1;
			P[16]=schimba;
			end
	
		2'b01:begin	
			P[16:0]=P+A;
			schimba=P[16];
			P=P>>1;
			P[16]=schimba;
			end
	
		2'b10:begin
			P[16:0]=P+S;
			schimba=P[16];
			P=P>>1;
			P[16]=schimba;
			end
			
		endcase	
	end
end	
	assign product=P[16:1];
endmodule	
	